module mos6502s_instruction_decoder(
  input [7:0] opcode,
  output [3:0] addr_mode,
  output [3:0] alu_op,
  output [3:0] instr_type,
  output [1:0] src_reg,
  output [1:0] dst_reg,
  output [2:0] branch_cond,
  output [2:0] cycles_base,
  output is_read,
  output is_write,
  output is_rmw,
  output sets_nz,
  output sets_c,
  output sets_v,
  output writes_reg,
  output is_status_op,
  output illegal
);

  assign addr_mode = ((opcode == 8'd105) ? 2'd2 : ((opcode == 8'd101) ? 2'd3 : ((opcode == 8'd117) ? 3'd4 : ((opcode == 8'd109) ? 3'd6 : ((opcode == 8'd125) ? 3'd7 : ((opcode == 8'd121) ? 4'd8 : ((opcode == 8'd97) ? 4'd10 : ((opcode == 8'd113) ? 4'd11 : ((opcode == 8'd233) ? 2'd2 : ((opcode == 8'd229) ? 2'd3 : ((opcode == 8'd245) ? 3'd4 : ((opcode == 8'd237) ? 3'd6 : ((opcode == 8'd253) ? 3'd7 : ((opcode == 8'd249) ? 4'd8 : ((opcode == 8'd225) ? 4'd10 : ((opcode == 8'd241) ? 4'd11 : ((opcode == 8'd41) ? 2'd2 : ((opcode == 8'd37) ? 2'd3 : ((opcode == 8'd53) ? 3'd4 : ((opcode == 8'd45) ? 3'd6 : ((opcode == 8'd61) ? 3'd7 : ((opcode == 8'd57) ? 4'd8 : ((opcode == 8'd33) ? 4'd10 : ((opcode == 8'd49) ? 4'd11 : ((opcode == 8'd9) ? 2'd2 : ((opcode == 8'd5) ? 2'd3 : ((opcode == 8'd21) ? 3'd4 : ((opcode == 8'd13) ? 3'd6 : ((opcode == 8'd29) ? 3'd7 : ((opcode == 8'd25) ? 4'd8 : ((opcode == 8'd1) ? 4'd10 : ((opcode == 8'd17) ? 4'd11 : ((opcode == 8'd73) ? 2'd2 : ((opcode == 8'd69) ? 2'd3 : ((opcode == 8'd85) ? 3'd4 : ((opcode == 8'd77) ? 3'd6 : ((opcode == 8'd93) ? 3'd7 : ((opcode == 8'd89) ? 4'd8 : ((opcode == 8'd65) ? 4'd10 : ((opcode == 8'd81) ? 4'd11 : ((opcode == 8'd201) ? 2'd2 : ((opcode == 8'd197) ? 2'd3 : ((opcode == 8'd213) ? 3'd4 : ((opcode == 8'd205) ? 3'd6 : ((opcode == 8'd221) ? 3'd7 : ((opcode == 8'd217) ? 4'd8 : ((opcode == 8'd193) ? 4'd10 : ((opcode == 8'd209) ? 4'd11 : ((opcode == 8'd224) ? 2'd2 : ((opcode == 8'd228) ? 2'd3 : ((opcode == 8'd236) ? 3'd6 : ((opcode == 8'd192) ? 2'd2 : ((opcode == 8'd196) ? 2'd3 : ((opcode == 8'd204) ? 3'd6 : ((opcode == 8'd36) ? 2'd3 : ((opcode == 8'd44) ? 3'd6 : ((opcode == 8'd169) ? 2'd2 : ((opcode == 8'd165) ? 2'd3 : ((opcode == 8'd181) ? 3'd4 : ((opcode == 8'd173) ? 3'd6 : ((opcode == 8'd189) ? 3'd7 : ((opcode == 8'd185) ? 4'd8 : ((opcode == 8'd161) ? 4'd10 : ((opcode == 8'd177) ? 4'd11 : ((opcode == 8'd162) ? 2'd2 : ((opcode == 8'd166) ? 2'd3 : ((opcode == 8'd182) ? 3'd5 : ((opcode == 8'd174) ? 3'd6 : ((opcode == 8'd190) ? 4'd8 : ((opcode == 8'd160) ? 2'd2 : ((opcode == 8'd164) ? 2'd3 : ((opcode == 8'd180) ? 3'd4 : ((opcode == 8'd172) ? 3'd6 : ((opcode == 8'd188) ? 3'd7 : ((opcode == 8'd133) ? 2'd3 : ((opcode == 8'd149) ? 3'd4 : ((opcode == 8'd141) ? 3'd6 : ((opcode == 8'd157) ? 3'd7 : ((opcode == 8'd153) ? 4'd8 : ((opcode == 8'd129) ? 4'd10 : ((opcode == 8'd145) ? 4'd11 : ((opcode == 8'd134) ? 2'd3 : ((opcode == 8'd150) ? 3'd5 : ((opcode == 8'd142) ? 3'd6 : ((opcode == 8'd132) ? 2'd3 : ((opcode == 8'd148) ? 3'd4 : ((opcode == 8'd140) ? 3'd6 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 2'd3 : ((opcode == 8'd246) ? 3'd4 : ((opcode == 8'd238) ? 3'd6 : ((opcode == 8'd254) ? 3'd7 : ((opcode == 8'd198) ? 2'd3 : ((opcode == 8'd214) ? 3'd4 : ((opcode == 8'd206) ? 3'd6 : ((opcode == 8'd222) ? 3'd7 : ((opcode == 8'd10) ? 1'b1 : ((opcode == 8'd6) ? 2'd3 : ((opcode == 8'd22) ? 3'd4 : ((opcode == 8'd14) ? 3'd6 : ((opcode == 8'd30) ? 3'd7 : ((opcode == 8'd74) ? 1'b1 : ((opcode == 8'd70) ? 2'd3 : ((opcode == 8'd86) ? 3'd4 : ((opcode == 8'd78) ? 3'd6 : ((opcode == 8'd94) ? 3'd7 : ((opcode == 8'd42) ? 1'b1 : ((opcode == 8'd38) ? 2'd3 : ((opcode == 8'd54) ? 3'd4 : ((opcode == 8'd46) ? 3'd6 : ((opcode == 8'd62) ? 3'd7 : ((opcode == 8'd106) ? 1'b1 : ((opcode == 8'd102) ? 2'd3 : ((opcode == 8'd118) ? 3'd4 : ((opcode == 8'd110) ? 3'd6 : ((opcode == 8'd126) ? 3'd7 : ((opcode == 8'd16) ? 4'd12 : ((opcode == 8'd48) ? 4'd12 : ((opcode == 8'd80) ? 4'd12 : ((opcode == 8'd112) ? 4'd12 : ((opcode == 8'd144) ? 4'd12 : ((opcode == 8'd176) ? 4'd12 : ((opcode == 8'd208) ? 4'd12 : ((opcode == 8'd240) ? 4'd12 : ((opcode == 8'd76) ? 3'd6 : ((opcode == 8'd108) ? 4'd9 : ((opcode == 8'd32) ? 3'd6 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign alu_op = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b1 : ((opcode == 8'd229) ? 1'b1 : ((opcode == 8'd245) ? 1'b1 : ((opcode == 8'd237) ? 1'b1 : ((opcode == 8'd253) ? 1'b1 : ((opcode == 8'd249) ? 1'b1 : ((opcode == 8'd225) ? 1'b1 : ((opcode == 8'd241) ? 1'b1 : ((opcode == 8'd41) ? 2'd2 : ((opcode == 8'd37) ? 2'd2 : ((opcode == 8'd53) ? 2'd2 : ((opcode == 8'd45) ? 2'd2 : ((opcode == 8'd61) ? 2'd2 : ((opcode == 8'd57) ? 2'd2 : ((opcode == 8'd33) ? 2'd2 : ((opcode == 8'd49) ? 2'd2 : ((opcode == 8'd9) ? 2'd3 : ((opcode == 8'd5) ? 2'd3 : ((opcode == 8'd21) ? 2'd3 : ((opcode == 8'd13) ? 2'd3 : ((opcode == 8'd29) ? 2'd3 : ((opcode == 8'd25) ? 2'd3 : ((opcode == 8'd1) ? 2'd3 : ((opcode == 8'd17) ? 2'd3 : ((opcode == 8'd73) ? 3'd4 : ((opcode == 8'd69) ? 3'd4 : ((opcode == 8'd85) ? 3'd4 : ((opcode == 8'd77) ? 3'd4 : ((opcode == 8'd93) ? 3'd4 : ((opcode == 8'd89) ? 3'd4 : ((opcode == 8'd65) ? 3'd4 : ((opcode == 8'd81) ? 3'd4 : ((opcode == 8'd201) ? 4'd11 : ((opcode == 8'd197) ? 4'd11 : ((opcode == 8'd213) ? 4'd11 : ((opcode == 8'd205) ? 4'd11 : ((opcode == 8'd221) ? 4'd11 : ((opcode == 8'd217) ? 4'd11 : ((opcode == 8'd193) ? 4'd11 : ((opcode == 8'd209) ? 4'd11 : ((opcode == 8'd224) ? 4'd11 : ((opcode == 8'd228) ? 4'd11 : ((opcode == 8'd236) ? 4'd11 : ((opcode == 8'd192) ? 4'd11 : ((opcode == 8'd196) ? 4'd11 : ((opcode == 8'd204) ? 4'd11 : ((opcode == 8'd36) ? 4'd12 : ((opcode == 8'd44) ? 4'd12 : ((opcode == 8'd169) ? 4'd13 : ((opcode == 8'd165) ? 4'd13 : ((opcode == 8'd181) ? 4'd13 : ((opcode == 8'd173) ? 4'd13 : ((opcode == 8'd189) ? 4'd13 : ((opcode == 8'd185) ? 4'd13 : ((opcode == 8'd161) ? 4'd13 : ((opcode == 8'd177) ? 4'd13 : ((opcode == 8'd162) ? 4'd13 : ((opcode == 8'd166) ? 4'd13 : ((opcode == 8'd182) ? 4'd13 : ((opcode == 8'd174) ? 4'd13 : ((opcode == 8'd190) ? 4'd13 : ((opcode == 8'd160) ? 4'd13 : ((opcode == 8'd164) ? 4'd13 : ((opcode == 8'd180) ? 4'd13 : ((opcode == 8'd172) ? 4'd13 : ((opcode == 8'd188) ? 4'd13 : ((opcode == 8'd133) ? 4'd15 : ((opcode == 8'd149) ? 4'd15 : ((opcode == 8'd141) ? 4'd15 : ((opcode == 8'd157) ? 4'd15 : ((opcode == 8'd153) ? 4'd15 : ((opcode == 8'd129) ? 4'd15 : ((opcode == 8'd145) ? 4'd15 : ((opcode == 8'd134) ? 4'd15 : ((opcode == 8'd150) ? 4'd15 : ((opcode == 8'd142) ? 4'd15 : ((opcode == 8'd132) ? 4'd15 : ((opcode == 8'd148) ? 4'd15 : ((opcode == 8'd140) ? 4'd15 : ((opcode == 8'd170) ? 4'd13 : ((opcode == 8'd138) ? 4'd13 : ((opcode == 8'd168) ? 4'd13 : ((opcode == 8'd152) ? 4'd13 : ((opcode == 8'd186) ? 4'd13 : ((opcode == 8'd154) ? 4'd13 : ((opcode == 8'd232) ? 4'd9 : ((opcode == 8'd202) ? 4'd10 : ((opcode == 8'd200) ? 4'd9 : ((opcode == 8'd136) ? 4'd10 : ((opcode == 8'd230) ? 4'd9 : ((opcode == 8'd246) ? 4'd9 : ((opcode == 8'd238) ? 4'd9 : ((opcode == 8'd254) ? 4'd9 : ((opcode == 8'd198) ? 4'd10 : ((opcode == 8'd214) ? 4'd10 : ((opcode == 8'd206) ? 4'd10 : ((opcode == 8'd222) ? 4'd10 : ((opcode == 8'd10) ? 3'd5 : ((opcode == 8'd6) ? 3'd5 : ((opcode == 8'd22) ? 3'd5 : ((opcode == 8'd14) ? 3'd5 : ((opcode == 8'd30) ? 3'd5 : ((opcode == 8'd74) ? 3'd6 : ((opcode == 8'd70) ? 3'd6 : ((opcode == 8'd86) ? 3'd6 : ((opcode == 8'd78) ? 3'd6 : ((opcode == 8'd94) ? 3'd6 : ((opcode == 8'd42) ? 3'd7 : ((opcode == 8'd38) ? 3'd7 : ((opcode == 8'd54) ? 3'd7 : ((opcode == 8'd46) ? 3'd7 : ((opcode == 8'd62) ? 3'd7 : ((opcode == 8'd106) ? 4'd8 : ((opcode == 8'd102) ? 4'd8 : ((opcode == 8'd118) ? 4'd8 : ((opcode == 8'd110) ? 4'd8 : ((opcode == 8'd126) ? 4'd8 : ((opcode == 8'd16) ? 4'd15 : ((opcode == 8'd48) ? 4'd15 : ((opcode == 8'd80) ? 4'd15 : ((opcode == 8'd112) ? 4'd15 : ((opcode == 8'd144) ? 4'd15 : ((opcode == 8'd176) ? 4'd15 : ((opcode == 8'd208) ? 4'd15 : ((opcode == 8'd240) ? 4'd15 : ((opcode == 8'd76) ? 4'd15 : ((opcode == 8'd108) ? 4'd15 : ((opcode == 8'd32) ? 4'd15 : ((opcode == 8'd96) ? 4'd15 : ((opcode == 8'd64) ? 4'd15 : ((opcode == 8'd72) ? 4'd13 : ((opcode == 8'd8) ? 4'd13 : ((opcode == 8'd104) ? 4'd13 : ((opcode == 8'd40) ? 4'd13 : ((opcode == 8'd24) ? 4'd15 : ((opcode == 8'd56) ? 4'd15 : ((opcode == 8'd88) ? 4'd15 : ((opcode == 8'd120) ? 4'd15 : ((opcode == 8'd184) ? 4'd15 : ((opcode == 8'd216) ? 4'd15 : ((opcode == 8'd248) ? 4'd15 : ((opcode == 8'd234) ? 4'd15 : ((opcode == 8'd0) ? 4'd15 : 4'd15)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign instr_type = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b1 : ((opcode == 8'd165) ? 1'b1 : ((opcode == 8'd181) ? 1'b1 : ((opcode == 8'd173) ? 1'b1 : ((opcode == 8'd189) ? 1'b1 : ((opcode == 8'd185) ? 1'b1 : ((opcode == 8'd161) ? 1'b1 : ((opcode == 8'd177) ? 1'b1 : ((opcode == 8'd162) ? 1'b1 : ((opcode == 8'd166) ? 1'b1 : ((opcode == 8'd182) ? 1'b1 : ((opcode == 8'd174) ? 1'b1 : ((opcode == 8'd190) ? 1'b1 : ((opcode == 8'd160) ? 1'b1 : ((opcode == 8'd164) ? 1'b1 : ((opcode == 8'd180) ? 1'b1 : ((opcode == 8'd172) ? 1'b1 : ((opcode == 8'd188) ? 1'b1 : ((opcode == 8'd133) ? 2'd2 : ((opcode == 8'd149) ? 2'd2 : ((opcode == 8'd141) ? 2'd2 : ((opcode == 8'd157) ? 2'd2 : ((opcode == 8'd153) ? 2'd2 : ((opcode == 8'd129) ? 2'd2 : ((opcode == 8'd145) ? 2'd2 : ((opcode == 8'd134) ? 2'd2 : ((opcode == 8'd150) ? 2'd2 : ((opcode == 8'd142) ? 2'd2 : ((opcode == 8'd132) ? 2'd2 : ((opcode == 8'd148) ? 2'd2 : ((opcode == 8'd140) ? 2'd2 : ((opcode == 8'd170) ? 2'd3 : ((opcode == 8'd138) ? 2'd3 : ((opcode == 8'd168) ? 2'd3 : ((opcode == 8'd152) ? 2'd3 : ((opcode == 8'd186) ? 2'd3 : ((opcode == 8'd154) ? 2'd3 : ((opcode == 8'd232) ? 3'd4 : ((opcode == 8'd202) ? 3'd4 : ((opcode == 8'd200) ? 3'd4 : ((opcode == 8'd136) ? 3'd4 : ((opcode == 8'd230) ? 3'd4 : ((opcode == 8'd246) ? 3'd4 : ((opcode == 8'd238) ? 3'd4 : ((opcode == 8'd254) ? 3'd4 : ((opcode == 8'd198) ? 3'd4 : ((opcode == 8'd214) ? 3'd4 : ((opcode == 8'd206) ? 3'd4 : ((opcode == 8'd222) ? 3'd4 : ((opcode == 8'd10) ? 3'd5 : ((opcode == 8'd6) ? 3'd5 : ((opcode == 8'd22) ? 3'd5 : ((opcode == 8'd14) ? 3'd5 : ((opcode == 8'd30) ? 3'd5 : ((opcode == 8'd74) ? 3'd5 : ((opcode == 8'd70) ? 3'd5 : ((opcode == 8'd86) ? 3'd5 : ((opcode == 8'd78) ? 3'd5 : ((opcode == 8'd94) ? 3'd5 : ((opcode == 8'd42) ? 3'd5 : ((opcode == 8'd38) ? 3'd5 : ((opcode == 8'd54) ? 3'd5 : ((opcode == 8'd46) ? 3'd5 : ((opcode == 8'd62) ? 3'd5 : ((opcode == 8'd106) ? 3'd5 : ((opcode == 8'd102) ? 3'd5 : ((opcode == 8'd118) ? 3'd5 : ((opcode == 8'd110) ? 3'd5 : ((opcode == 8'd126) ? 3'd5 : ((opcode == 8'd16) ? 3'd6 : ((opcode == 8'd48) ? 3'd6 : ((opcode == 8'd80) ? 3'd6 : ((opcode == 8'd112) ? 3'd6 : ((opcode == 8'd144) ? 3'd6 : ((opcode == 8'd176) ? 3'd6 : ((opcode == 8'd208) ? 3'd6 : ((opcode == 8'd240) ? 3'd6 : ((opcode == 8'd76) ? 3'd7 : ((opcode == 8'd108) ? 3'd7 : ((opcode == 8'd32) ? 3'd7 : ((opcode == 8'd96) ? 3'd7 : ((opcode == 8'd64) ? 3'd7 : ((opcode == 8'd72) ? 4'd8 : ((opcode == 8'd8) ? 4'd8 : ((opcode == 8'd104) ? 4'd8 : ((opcode == 8'd40) ? 4'd8 : ((opcode == 8'd24) ? 4'd9 : ((opcode == 8'd56) ? 4'd9 : ((opcode == 8'd88) ? 4'd9 : ((opcode == 8'd120) ? 4'd9 : ((opcode == 8'd184) ? 4'd9 : ((opcode == 8'd216) ? 4'd9 : ((opcode == 8'd248) ? 4'd9 : ((opcode == 8'd234) ? 4'd10 : ((opcode == 8'd0) ? 4'd11 : 4'd10)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign src_reg = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b1 : ((opcode == 8'd228) ? 1'b1 : ((opcode == 8'd236) ? 1'b1 : ((opcode == 8'd192) ? 2'd2 : ((opcode == 8'd196) ? 2'd2 : ((opcode == 8'd204) ? 2'd2 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b1 : ((opcode == 8'd166) ? 1'b1 : ((opcode == 8'd182) ? 1'b1 : ((opcode == 8'd174) ? 1'b1 : ((opcode == 8'd190) ? 1'b1 : ((opcode == 8'd160) ? 2'd2 : ((opcode == 8'd164) ? 2'd2 : ((opcode == 8'd180) ? 2'd2 : ((opcode == 8'd172) ? 2'd2 : ((opcode == 8'd188) ? 2'd2 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b1 : ((opcode == 8'd150) ? 1'b1 : ((opcode == 8'd142) ? 1'b1 : ((opcode == 8'd132) ? 2'd2 : ((opcode == 8'd148) ? 2'd2 : ((opcode == 8'd140) ? 2'd2 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b1 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 2'd2 : ((opcode == 8'd186) ? 1'b1 : ((opcode == 8'd154) ? 1'b1 : ((opcode == 8'd232) ? 1'b1 : ((opcode == 8'd202) ? 1'b1 : ((opcode == 8'd200) ? 2'd2 : ((opcode == 8'd136) ? 2'd2 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign dst_reg = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b1 : ((opcode == 8'd228) ? 1'b1 : ((opcode == 8'd236) ? 1'b1 : ((opcode == 8'd192) ? 2'd2 : ((opcode == 8'd196) ? 2'd2 : ((opcode == 8'd204) ? 2'd2 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b1 : ((opcode == 8'd166) ? 1'b1 : ((opcode == 8'd182) ? 1'b1 : ((opcode == 8'd174) ? 1'b1 : ((opcode == 8'd190) ? 1'b1 : ((opcode == 8'd160) ? 2'd2 : ((opcode == 8'd164) ? 2'd2 : ((opcode == 8'd180) ? 2'd2 : ((opcode == 8'd172) ? 2'd2 : ((opcode == 8'd188) ? 2'd2 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b1 : ((opcode == 8'd150) ? 1'b1 : ((opcode == 8'd142) ? 1'b1 : ((opcode == 8'd132) ? 2'd2 : ((opcode == 8'd148) ? 2'd2 : ((opcode == 8'd140) ? 2'd2 : ((opcode == 8'd170) ? 1'b1 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 2'd2 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b1 : ((opcode == 8'd154) ? 1'b1 : ((opcode == 8'd232) ? 1'b1 : ((opcode == 8'd202) ? 1'b1 : ((opcode == 8'd200) ? 2'd2 : ((opcode == 8'd136) ? 2'd2 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign branch_cond = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b1 : ((opcode == 8'd80) ? 2'd2 : ((opcode == 8'd112) ? 2'd3 : ((opcode == 8'd144) ? 3'd4 : ((opcode == 8'd176) ? 3'd5 : ((opcode == 8'd208) ? 3'd6 : ((opcode == 8'd240) ? 3'd7 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign cycles_base = ((opcode == 8'd105) ? 2'd2 : ((opcode == 8'd101) ? 2'd3 : ((opcode == 8'd117) ? 3'd4 : ((opcode == 8'd109) ? 3'd4 : ((opcode == 8'd125) ? 3'd4 : ((opcode == 8'd121) ? 3'd4 : ((opcode == 8'd97) ? 3'd6 : ((opcode == 8'd113) ? 3'd5 : ((opcode == 8'd233) ? 2'd2 : ((opcode == 8'd229) ? 2'd3 : ((opcode == 8'd245) ? 3'd4 : ((opcode == 8'd237) ? 3'd4 : ((opcode == 8'd253) ? 3'd4 : ((opcode == 8'd249) ? 3'd4 : ((opcode == 8'd225) ? 3'd6 : ((opcode == 8'd241) ? 3'd5 : ((opcode == 8'd41) ? 2'd2 : ((opcode == 8'd37) ? 2'd3 : ((opcode == 8'd53) ? 3'd4 : ((opcode == 8'd45) ? 3'd4 : ((opcode == 8'd61) ? 3'd4 : ((opcode == 8'd57) ? 3'd4 : ((opcode == 8'd33) ? 3'd6 : ((opcode == 8'd49) ? 3'd5 : ((opcode == 8'd9) ? 2'd2 : ((opcode == 8'd5) ? 2'd3 : ((opcode == 8'd21) ? 3'd4 : ((opcode == 8'd13) ? 3'd4 : ((opcode == 8'd29) ? 3'd4 : ((opcode == 8'd25) ? 3'd4 : ((opcode == 8'd1) ? 3'd6 : ((opcode == 8'd17) ? 3'd5 : ((opcode == 8'd73) ? 2'd2 : ((opcode == 8'd69) ? 2'd3 : ((opcode == 8'd85) ? 3'd4 : ((opcode == 8'd77) ? 3'd4 : ((opcode == 8'd93) ? 3'd4 : ((opcode == 8'd89) ? 3'd4 : ((opcode == 8'd65) ? 3'd6 : ((opcode == 8'd81) ? 3'd5 : ((opcode == 8'd201) ? 2'd2 : ((opcode == 8'd197) ? 2'd3 : ((opcode == 8'd213) ? 3'd4 : ((opcode == 8'd205) ? 3'd4 : ((opcode == 8'd221) ? 3'd4 : ((opcode == 8'd217) ? 3'd4 : ((opcode == 8'd193) ? 3'd6 : ((opcode == 8'd209) ? 3'd5 : ((opcode == 8'd224) ? 2'd2 : ((opcode == 8'd228) ? 2'd3 : ((opcode == 8'd236) ? 3'd4 : ((opcode == 8'd192) ? 2'd2 : ((opcode == 8'd196) ? 2'd3 : ((opcode == 8'd204) ? 3'd4 : ((opcode == 8'd36) ? 2'd3 : ((opcode == 8'd44) ? 3'd4 : ((opcode == 8'd169) ? 2'd2 : ((opcode == 8'd165) ? 2'd3 : ((opcode == 8'd181) ? 3'd4 : ((opcode == 8'd173) ? 3'd4 : ((opcode == 8'd189) ? 3'd4 : ((opcode == 8'd185) ? 3'd4 : ((opcode == 8'd161) ? 3'd6 : ((opcode == 8'd177) ? 3'd5 : ((opcode == 8'd162) ? 2'd2 : ((opcode == 8'd166) ? 2'd3 : ((opcode == 8'd182) ? 3'd4 : ((opcode == 8'd174) ? 3'd4 : ((opcode == 8'd190) ? 3'd4 : ((opcode == 8'd160) ? 2'd2 : ((opcode == 8'd164) ? 2'd3 : ((opcode == 8'd180) ? 3'd4 : ((opcode == 8'd172) ? 3'd4 : ((opcode == 8'd188) ? 3'd4 : ((opcode == 8'd133) ? 2'd3 : ((opcode == 8'd149) ? 3'd4 : ((opcode == 8'd141) ? 3'd4 : ((opcode == 8'd157) ? 3'd5 : ((opcode == 8'd153) ? 3'd5 : ((opcode == 8'd129) ? 3'd6 : ((opcode == 8'd145) ? 3'd6 : ((opcode == 8'd134) ? 2'd3 : ((opcode == 8'd150) ? 3'd4 : ((opcode == 8'd142) ? 3'd4 : ((opcode == 8'd132) ? 2'd3 : ((opcode == 8'd148) ? 3'd4 : ((opcode == 8'd140) ? 3'd4 : ((opcode == 8'd170) ? 2'd2 : ((opcode == 8'd138) ? 2'd2 : ((opcode == 8'd168) ? 2'd2 : ((opcode == 8'd152) ? 2'd2 : ((opcode == 8'd186) ? 2'd2 : ((opcode == 8'd154) ? 2'd2 : ((opcode == 8'd232) ? 2'd2 : ((opcode == 8'd202) ? 2'd2 : ((opcode == 8'd200) ? 2'd2 : ((opcode == 8'd136) ? 2'd2 : ((opcode == 8'd230) ? 3'd5 : ((opcode == 8'd246) ? 3'd6 : ((opcode == 8'd238) ? 3'd6 : ((opcode == 8'd254) ? 3'd7 : ((opcode == 8'd198) ? 3'd5 : ((opcode == 8'd214) ? 3'd6 : ((opcode == 8'd206) ? 3'd6 : ((opcode == 8'd222) ? 3'd7 : ((opcode == 8'd10) ? 2'd2 : ((opcode == 8'd6) ? 3'd5 : ((opcode == 8'd22) ? 3'd6 : ((opcode == 8'd14) ? 3'd6 : ((opcode == 8'd30) ? 3'd7 : ((opcode == 8'd74) ? 2'd2 : ((opcode == 8'd70) ? 3'd5 : ((opcode == 8'd86) ? 3'd6 : ((opcode == 8'd78) ? 3'd6 : ((opcode == 8'd94) ? 3'd7 : ((opcode == 8'd42) ? 2'd2 : ((opcode == 8'd38) ? 3'd5 : ((opcode == 8'd54) ? 3'd6 : ((opcode == 8'd46) ? 3'd6 : ((opcode == 8'd62) ? 3'd7 : ((opcode == 8'd106) ? 2'd2 : ((opcode == 8'd102) ? 3'd5 : ((opcode == 8'd118) ? 3'd6 : ((opcode == 8'd110) ? 3'd6 : ((opcode == 8'd126) ? 3'd7 : ((opcode == 8'd16) ? 2'd2 : ((opcode == 8'd48) ? 2'd2 : ((opcode == 8'd80) ? 2'd2 : ((opcode == 8'd112) ? 2'd2 : ((opcode == 8'd144) ? 2'd2 : ((opcode == 8'd176) ? 2'd2 : ((opcode == 8'd208) ? 2'd2 : ((opcode == 8'd240) ? 2'd2 : ((opcode == 8'd76) ? 2'd3 : ((opcode == 8'd108) ? 3'd5 : ((opcode == 8'd32) ? 3'd6 : ((opcode == 8'd96) ? 3'd6 : ((opcode == 8'd64) ? 3'd6 : ((opcode == 8'd72) ? 2'd3 : ((opcode == 8'd8) ? 2'd3 : ((opcode == 8'd104) ? 3'd4 : ((opcode == 8'd40) ? 3'd4 : ((opcode == 8'd24) ? 2'd2 : ((opcode == 8'd56) ? 2'd2 : ((opcode == 8'd88) ? 2'd2 : ((opcode == 8'd120) ? 2'd2 : ((opcode == 8'd184) ? 2'd2 : ((opcode == 8'd216) ? 2'd2 : ((opcode == 8'd248) ? 2'd2 : ((opcode == 8'd234) ? 2'd2 : ((opcode == 8'd0) ? 3'd7 : 2'd2)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign is_read = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b1 : ((opcode == 8'd117) ? 1'b1 : ((opcode == 8'd109) ? 1'b1 : ((opcode == 8'd125) ? 1'b1 : ((opcode == 8'd121) ? 1'b1 : ((opcode == 8'd97) ? 1'b1 : ((opcode == 8'd113) ? 1'b1 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b1 : ((opcode == 8'd245) ? 1'b1 : ((opcode == 8'd237) ? 1'b1 : ((opcode == 8'd253) ? 1'b1 : ((opcode == 8'd249) ? 1'b1 : ((opcode == 8'd225) ? 1'b1 : ((opcode == 8'd241) ? 1'b1 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b1 : ((opcode == 8'd53) ? 1'b1 : ((opcode == 8'd45) ? 1'b1 : ((opcode == 8'd61) ? 1'b1 : ((opcode == 8'd57) ? 1'b1 : ((opcode == 8'd33) ? 1'b1 : ((opcode == 8'd49) ? 1'b1 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b1 : ((opcode == 8'd21) ? 1'b1 : ((opcode == 8'd13) ? 1'b1 : ((opcode == 8'd29) ? 1'b1 : ((opcode == 8'd25) ? 1'b1 : ((opcode == 8'd1) ? 1'b1 : ((opcode == 8'd17) ? 1'b1 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b1 : ((opcode == 8'd85) ? 1'b1 : ((opcode == 8'd77) ? 1'b1 : ((opcode == 8'd93) ? 1'b1 : ((opcode == 8'd89) ? 1'b1 : ((opcode == 8'd65) ? 1'b1 : ((opcode == 8'd81) ? 1'b1 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b1 : ((opcode == 8'd213) ? 1'b1 : ((opcode == 8'd205) ? 1'b1 : ((opcode == 8'd221) ? 1'b1 : ((opcode == 8'd217) ? 1'b1 : ((opcode == 8'd193) ? 1'b1 : ((opcode == 8'd209) ? 1'b1 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b1 : ((opcode == 8'd236) ? 1'b1 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b1 : ((opcode == 8'd204) ? 1'b1 : ((opcode == 8'd36) ? 1'b1 : ((opcode == 8'd44) ? 1'b1 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b1 : ((opcode == 8'd181) ? 1'b1 : ((opcode == 8'd173) ? 1'b1 : ((opcode == 8'd189) ? 1'b1 : ((opcode == 8'd185) ? 1'b1 : ((opcode == 8'd161) ? 1'b1 : ((opcode == 8'd177) ? 1'b1 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b1 : ((opcode == 8'd182) ? 1'b1 : ((opcode == 8'd174) ? 1'b1 : ((opcode == 8'd190) ? 1'b1 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b1 : ((opcode == 8'd180) ? 1'b1 : ((opcode == 8'd172) ? 1'b1 : ((opcode == 8'd188) ? 1'b1 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b1 : ((opcode == 8'd246) ? 1'b1 : ((opcode == 8'd238) ? 1'b1 : ((opcode == 8'd254) ? 1'b1 : ((opcode == 8'd198) ? 1'b1 : ((opcode == 8'd214) ? 1'b1 : ((opcode == 8'd206) ? 1'b1 : ((opcode == 8'd222) ? 1'b1 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b1 : ((opcode == 8'd22) ? 1'b1 : ((opcode == 8'd14) ? 1'b1 : ((opcode == 8'd30) ? 1'b1 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b1 : ((opcode == 8'd86) ? 1'b1 : ((opcode == 8'd78) ? 1'b1 : ((opcode == 8'd94) ? 1'b1 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b1 : ((opcode == 8'd54) ? 1'b1 : ((opcode == 8'd46) ? 1'b1 : ((opcode == 8'd62) ? 1'b1 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b1 : ((opcode == 8'd118) ? 1'b1 : ((opcode == 8'd110) ? 1'b1 : ((opcode == 8'd126) ? 1'b1 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b1 : ((opcode == 8'd40) ? 1'b1 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign is_write = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b1 : ((opcode == 8'd149) ? 1'b1 : ((opcode == 8'd141) ? 1'b1 : ((opcode == 8'd157) ? 1'b1 : ((opcode == 8'd153) ? 1'b1 : ((opcode == 8'd129) ? 1'b1 : ((opcode == 8'd145) ? 1'b1 : ((opcode == 8'd134) ? 1'b1 : ((opcode == 8'd150) ? 1'b1 : ((opcode == 8'd142) ? 1'b1 : ((opcode == 8'd132) ? 1'b1 : ((opcode == 8'd148) ? 1'b1 : ((opcode == 8'd140) ? 1'b1 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b1 : ((opcode == 8'd246) ? 1'b1 : ((opcode == 8'd238) ? 1'b1 : ((opcode == 8'd254) ? 1'b1 : ((opcode == 8'd198) ? 1'b1 : ((opcode == 8'd214) ? 1'b1 : ((opcode == 8'd206) ? 1'b1 : ((opcode == 8'd222) ? 1'b1 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b1 : ((opcode == 8'd22) ? 1'b1 : ((opcode == 8'd14) ? 1'b1 : ((opcode == 8'd30) ? 1'b1 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b1 : ((opcode == 8'd86) ? 1'b1 : ((opcode == 8'd78) ? 1'b1 : ((opcode == 8'd94) ? 1'b1 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b1 : ((opcode == 8'd54) ? 1'b1 : ((opcode == 8'd46) ? 1'b1 : ((opcode == 8'd62) ? 1'b1 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b1 : ((opcode == 8'd118) ? 1'b1 : ((opcode == 8'd110) ? 1'b1 : ((opcode == 8'd126) ? 1'b1 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b1 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b1 : ((opcode == 8'd8) ? 1'b1 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign is_rmw = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b1 : ((opcode == 8'd246) ? 1'b1 : ((opcode == 8'd238) ? 1'b1 : ((opcode == 8'd254) ? 1'b1 : ((opcode == 8'd198) ? 1'b1 : ((opcode == 8'd214) ? 1'b1 : ((opcode == 8'd206) ? 1'b1 : ((opcode == 8'd222) ? 1'b1 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b1 : ((opcode == 8'd22) ? 1'b1 : ((opcode == 8'd14) ? 1'b1 : ((opcode == 8'd30) ? 1'b1 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b1 : ((opcode == 8'd86) ? 1'b1 : ((opcode == 8'd78) ? 1'b1 : ((opcode == 8'd94) ? 1'b1 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b1 : ((opcode == 8'd54) ? 1'b1 : ((opcode == 8'd46) ? 1'b1 : ((opcode == 8'd62) ? 1'b1 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b1 : ((opcode == 8'd118) ? 1'b1 : ((opcode == 8'd110) ? 1'b1 : ((opcode == 8'd126) ? 1'b1 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign sets_nz = ((opcode == 8'd105) ? 1'b1 : ((opcode == 8'd101) ? 1'b1 : ((opcode == 8'd117) ? 1'b1 : ((opcode == 8'd109) ? 1'b1 : ((opcode == 8'd125) ? 1'b1 : ((opcode == 8'd121) ? 1'b1 : ((opcode == 8'd97) ? 1'b1 : ((opcode == 8'd113) ? 1'b1 : ((opcode == 8'd233) ? 1'b1 : ((opcode == 8'd229) ? 1'b1 : ((opcode == 8'd245) ? 1'b1 : ((opcode == 8'd237) ? 1'b1 : ((opcode == 8'd253) ? 1'b1 : ((opcode == 8'd249) ? 1'b1 : ((opcode == 8'd225) ? 1'b1 : ((opcode == 8'd241) ? 1'b1 : ((opcode == 8'd41) ? 1'b1 : ((opcode == 8'd37) ? 1'b1 : ((opcode == 8'd53) ? 1'b1 : ((opcode == 8'd45) ? 1'b1 : ((opcode == 8'd61) ? 1'b1 : ((opcode == 8'd57) ? 1'b1 : ((opcode == 8'd33) ? 1'b1 : ((opcode == 8'd49) ? 1'b1 : ((opcode == 8'd9) ? 1'b1 : ((opcode == 8'd5) ? 1'b1 : ((opcode == 8'd21) ? 1'b1 : ((opcode == 8'd13) ? 1'b1 : ((opcode == 8'd29) ? 1'b1 : ((opcode == 8'd25) ? 1'b1 : ((opcode == 8'd1) ? 1'b1 : ((opcode == 8'd17) ? 1'b1 : ((opcode == 8'd73) ? 1'b1 : ((opcode == 8'd69) ? 1'b1 : ((opcode == 8'd85) ? 1'b1 : ((opcode == 8'd77) ? 1'b1 : ((opcode == 8'd93) ? 1'b1 : ((opcode == 8'd89) ? 1'b1 : ((opcode == 8'd65) ? 1'b1 : ((opcode == 8'd81) ? 1'b1 : ((opcode == 8'd201) ? 1'b1 : ((opcode == 8'd197) ? 1'b1 : ((opcode == 8'd213) ? 1'b1 : ((opcode == 8'd205) ? 1'b1 : ((opcode == 8'd221) ? 1'b1 : ((opcode == 8'd217) ? 1'b1 : ((opcode == 8'd193) ? 1'b1 : ((opcode == 8'd209) ? 1'b1 : ((opcode == 8'd224) ? 1'b1 : ((opcode == 8'd228) ? 1'b1 : ((opcode == 8'd236) ? 1'b1 : ((opcode == 8'd192) ? 1'b1 : ((opcode == 8'd196) ? 1'b1 : ((opcode == 8'd204) ? 1'b1 : ((opcode == 8'd36) ? 1'b1 : ((opcode == 8'd44) ? 1'b1 : ((opcode == 8'd169) ? 1'b1 : ((opcode == 8'd165) ? 1'b1 : ((opcode == 8'd181) ? 1'b1 : ((opcode == 8'd173) ? 1'b1 : ((opcode == 8'd189) ? 1'b1 : ((opcode == 8'd185) ? 1'b1 : ((opcode == 8'd161) ? 1'b1 : ((opcode == 8'd177) ? 1'b1 : ((opcode == 8'd162) ? 1'b1 : ((opcode == 8'd166) ? 1'b1 : ((opcode == 8'd182) ? 1'b1 : ((opcode == 8'd174) ? 1'b1 : ((opcode == 8'd190) ? 1'b1 : ((opcode == 8'd160) ? 1'b1 : ((opcode == 8'd164) ? 1'b1 : ((opcode == 8'd180) ? 1'b1 : ((opcode == 8'd172) ? 1'b1 : ((opcode == 8'd188) ? 1'b1 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b1 : ((opcode == 8'd138) ? 1'b1 : ((opcode == 8'd168) ? 1'b1 : ((opcode == 8'd152) ? 1'b1 : ((opcode == 8'd186) ? 1'b1 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b1 : ((opcode == 8'd202) ? 1'b1 : ((opcode == 8'd200) ? 1'b1 : ((opcode == 8'd136) ? 1'b1 : ((opcode == 8'd230) ? 1'b1 : ((opcode == 8'd246) ? 1'b1 : ((opcode == 8'd238) ? 1'b1 : ((opcode == 8'd254) ? 1'b1 : ((opcode == 8'd198) ? 1'b1 : ((opcode == 8'd214) ? 1'b1 : ((opcode == 8'd206) ? 1'b1 : ((opcode == 8'd222) ? 1'b1 : ((opcode == 8'd10) ? 1'b1 : ((opcode == 8'd6) ? 1'b1 : ((opcode == 8'd22) ? 1'b1 : ((opcode == 8'd14) ? 1'b1 : ((opcode == 8'd30) ? 1'b1 : ((opcode == 8'd74) ? 1'b1 : ((opcode == 8'd70) ? 1'b1 : ((opcode == 8'd86) ? 1'b1 : ((opcode == 8'd78) ? 1'b1 : ((opcode == 8'd94) ? 1'b1 : ((opcode == 8'd42) ? 1'b1 : ((opcode == 8'd38) ? 1'b1 : ((opcode == 8'd54) ? 1'b1 : ((opcode == 8'd46) ? 1'b1 : ((opcode == 8'd62) ? 1'b1 : ((opcode == 8'd106) ? 1'b1 : ((opcode == 8'd102) ? 1'b1 : ((opcode == 8'd118) ? 1'b1 : ((opcode == 8'd110) ? 1'b1 : ((opcode == 8'd126) ? 1'b1 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b1 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign sets_c = ((opcode == 8'd105) ? 1'b1 : ((opcode == 8'd101) ? 1'b1 : ((opcode == 8'd117) ? 1'b1 : ((opcode == 8'd109) ? 1'b1 : ((opcode == 8'd125) ? 1'b1 : ((opcode == 8'd121) ? 1'b1 : ((opcode == 8'd97) ? 1'b1 : ((opcode == 8'd113) ? 1'b1 : ((opcode == 8'd233) ? 1'b1 : ((opcode == 8'd229) ? 1'b1 : ((opcode == 8'd245) ? 1'b1 : ((opcode == 8'd237) ? 1'b1 : ((opcode == 8'd253) ? 1'b1 : ((opcode == 8'd249) ? 1'b1 : ((opcode == 8'd225) ? 1'b1 : ((opcode == 8'd241) ? 1'b1 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b1 : ((opcode == 8'd197) ? 1'b1 : ((opcode == 8'd213) ? 1'b1 : ((opcode == 8'd205) ? 1'b1 : ((opcode == 8'd221) ? 1'b1 : ((opcode == 8'd217) ? 1'b1 : ((opcode == 8'd193) ? 1'b1 : ((opcode == 8'd209) ? 1'b1 : ((opcode == 8'd224) ? 1'b1 : ((opcode == 8'd228) ? 1'b1 : ((opcode == 8'd236) ? 1'b1 : ((opcode == 8'd192) ? 1'b1 : ((opcode == 8'd196) ? 1'b1 : ((opcode == 8'd204) ? 1'b1 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b1 : ((opcode == 8'd6) ? 1'b1 : ((opcode == 8'd22) ? 1'b1 : ((opcode == 8'd14) ? 1'b1 : ((opcode == 8'd30) ? 1'b1 : ((opcode == 8'd74) ? 1'b1 : ((opcode == 8'd70) ? 1'b1 : ((opcode == 8'd86) ? 1'b1 : ((opcode == 8'd78) ? 1'b1 : ((opcode == 8'd94) ? 1'b1 : ((opcode == 8'd42) ? 1'b1 : ((opcode == 8'd38) ? 1'b1 : ((opcode == 8'd54) ? 1'b1 : ((opcode == 8'd46) ? 1'b1 : ((opcode == 8'd62) ? 1'b1 : ((opcode == 8'd106) ? 1'b1 : ((opcode == 8'd102) ? 1'b1 : ((opcode == 8'd118) ? 1'b1 : ((opcode == 8'd110) ? 1'b1 : ((opcode == 8'd126) ? 1'b1 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b1 : ((opcode == 8'd24) ? 1'b1 : ((opcode == 8'd56) ? 1'b1 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign sets_v = ((opcode == 8'd105) ? 1'b1 : ((opcode == 8'd101) ? 1'b1 : ((opcode == 8'd117) ? 1'b1 : ((opcode == 8'd109) ? 1'b1 : ((opcode == 8'd125) ? 1'b1 : ((opcode == 8'd121) ? 1'b1 : ((opcode == 8'd97) ? 1'b1 : ((opcode == 8'd113) ? 1'b1 : ((opcode == 8'd233) ? 1'b1 : ((opcode == 8'd229) ? 1'b1 : ((opcode == 8'd245) ? 1'b1 : ((opcode == 8'd237) ? 1'b1 : ((opcode == 8'd253) ? 1'b1 : ((opcode == 8'd249) ? 1'b1 : ((opcode == 8'd225) ? 1'b1 : ((opcode == 8'd241) ? 1'b1 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b1 : ((opcode == 8'd44) ? 1'b1 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b1 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b1 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign writes_reg = ((opcode == 8'd105) ? 1'b1 : ((opcode == 8'd101) ? 1'b1 : ((opcode == 8'd117) ? 1'b1 : ((opcode == 8'd109) ? 1'b1 : ((opcode == 8'd125) ? 1'b1 : ((opcode == 8'd121) ? 1'b1 : ((opcode == 8'd97) ? 1'b1 : ((opcode == 8'd113) ? 1'b1 : ((opcode == 8'd233) ? 1'b1 : ((opcode == 8'd229) ? 1'b1 : ((opcode == 8'd245) ? 1'b1 : ((opcode == 8'd237) ? 1'b1 : ((opcode == 8'd253) ? 1'b1 : ((opcode == 8'd249) ? 1'b1 : ((opcode == 8'd225) ? 1'b1 : ((opcode == 8'd241) ? 1'b1 : ((opcode == 8'd41) ? 1'b1 : ((opcode == 8'd37) ? 1'b1 : ((opcode == 8'd53) ? 1'b1 : ((opcode == 8'd45) ? 1'b1 : ((opcode == 8'd61) ? 1'b1 : ((opcode == 8'd57) ? 1'b1 : ((opcode == 8'd33) ? 1'b1 : ((opcode == 8'd49) ? 1'b1 : ((opcode == 8'd9) ? 1'b1 : ((opcode == 8'd5) ? 1'b1 : ((opcode == 8'd21) ? 1'b1 : ((opcode == 8'd13) ? 1'b1 : ((opcode == 8'd29) ? 1'b1 : ((opcode == 8'd25) ? 1'b1 : ((opcode == 8'd1) ? 1'b1 : ((opcode == 8'd17) ? 1'b1 : ((opcode == 8'd73) ? 1'b1 : ((opcode == 8'd69) ? 1'b1 : ((opcode == 8'd85) ? 1'b1 : ((opcode == 8'd77) ? 1'b1 : ((opcode == 8'd93) ? 1'b1 : ((opcode == 8'd89) ? 1'b1 : ((opcode == 8'd65) ? 1'b1 : ((opcode == 8'd81) ? 1'b1 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b1 : ((opcode == 8'd165) ? 1'b1 : ((opcode == 8'd181) ? 1'b1 : ((opcode == 8'd173) ? 1'b1 : ((opcode == 8'd189) ? 1'b1 : ((opcode == 8'd185) ? 1'b1 : ((opcode == 8'd161) ? 1'b1 : ((opcode == 8'd177) ? 1'b1 : ((opcode == 8'd162) ? 1'b1 : ((opcode == 8'd166) ? 1'b1 : ((opcode == 8'd182) ? 1'b1 : ((opcode == 8'd174) ? 1'b1 : ((opcode == 8'd190) ? 1'b1 : ((opcode == 8'd160) ? 1'b1 : ((opcode == 8'd164) ? 1'b1 : ((opcode == 8'd180) ? 1'b1 : ((opcode == 8'd172) ? 1'b1 : ((opcode == 8'd188) ? 1'b1 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b1 : ((opcode == 8'd138) ? 1'b1 : ((opcode == 8'd168) ? 1'b1 : ((opcode == 8'd152) ? 1'b1 : ((opcode == 8'd186) ? 1'b1 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b1 : ((opcode == 8'd202) ? 1'b1 : ((opcode == 8'd200) ? 1'b1 : ((opcode == 8'd136) ? 1'b1 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b1 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b1 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b1 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b1 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b1 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign is_status_op = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b1 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b1 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
  assign illegal = ((opcode == 8'd105) ? 1'b0 : ((opcode == 8'd101) ? 1'b0 : ((opcode == 8'd117) ? 1'b0 : ((opcode == 8'd109) ? 1'b0 : ((opcode == 8'd125) ? 1'b0 : ((opcode == 8'd121) ? 1'b0 : ((opcode == 8'd97) ? 1'b0 : ((opcode == 8'd113) ? 1'b0 : ((opcode == 8'd233) ? 1'b0 : ((opcode == 8'd229) ? 1'b0 : ((opcode == 8'd245) ? 1'b0 : ((opcode == 8'd237) ? 1'b0 : ((opcode == 8'd253) ? 1'b0 : ((opcode == 8'd249) ? 1'b0 : ((opcode == 8'd225) ? 1'b0 : ((opcode == 8'd241) ? 1'b0 : ((opcode == 8'd41) ? 1'b0 : ((opcode == 8'd37) ? 1'b0 : ((opcode == 8'd53) ? 1'b0 : ((opcode == 8'd45) ? 1'b0 : ((opcode == 8'd61) ? 1'b0 : ((opcode == 8'd57) ? 1'b0 : ((opcode == 8'd33) ? 1'b0 : ((opcode == 8'd49) ? 1'b0 : ((opcode == 8'd9) ? 1'b0 : ((opcode == 8'd5) ? 1'b0 : ((opcode == 8'd21) ? 1'b0 : ((opcode == 8'd13) ? 1'b0 : ((opcode == 8'd29) ? 1'b0 : ((opcode == 8'd25) ? 1'b0 : ((opcode == 8'd1) ? 1'b0 : ((opcode == 8'd17) ? 1'b0 : ((opcode == 8'd73) ? 1'b0 : ((opcode == 8'd69) ? 1'b0 : ((opcode == 8'd85) ? 1'b0 : ((opcode == 8'd77) ? 1'b0 : ((opcode == 8'd93) ? 1'b0 : ((opcode == 8'd89) ? 1'b0 : ((opcode == 8'd65) ? 1'b0 : ((opcode == 8'd81) ? 1'b0 : ((opcode == 8'd201) ? 1'b0 : ((opcode == 8'd197) ? 1'b0 : ((opcode == 8'd213) ? 1'b0 : ((opcode == 8'd205) ? 1'b0 : ((opcode == 8'd221) ? 1'b0 : ((opcode == 8'd217) ? 1'b0 : ((opcode == 8'd193) ? 1'b0 : ((opcode == 8'd209) ? 1'b0 : ((opcode == 8'd224) ? 1'b0 : ((opcode == 8'd228) ? 1'b0 : ((opcode == 8'd236) ? 1'b0 : ((opcode == 8'd192) ? 1'b0 : ((opcode == 8'd196) ? 1'b0 : ((opcode == 8'd204) ? 1'b0 : ((opcode == 8'd36) ? 1'b0 : ((opcode == 8'd44) ? 1'b0 : ((opcode == 8'd169) ? 1'b0 : ((opcode == 8'd165) ? 1'b0 : ((opcode == 8'd181) ? 1'b0 : ((opcode == 8'd173) ? 1'b0 : ((opcode == 8'd189) ? 1'b0 : ((opcode == 8'd185) ? 1'b0 : ((opcode == 8'd161) ? 1'b0 : ((opcode == 8'd177) ? 1'b0 : ((opcode == 8'd162) ? 1'b0 : ((opcode == 8'd166) ? 1'b0 : ((opcode == 8'd182) ? 1'b0 : ((opcode == 8'd174) ? 1'b0 : ((opcode == 8'd190) ? 1'b0 : ((opcode == 8'd160) ? 1'b0 : ((opcode == 8'd164) ? 1'b0 : ((opcode == 8'd180) ? 1'b0 : ((opcode == 8'd172) ? 1'b0 : ((opcode == 8'd188) ? 1'b0 : ((opcode == 8'd133) ? 1'b0 : ((opcode == 8'd149) ? 1'b0 : ((opcode == 8'd141) ? 1'b0 : ((opcode == 8'd157) ? 1'b0 : ((opcode == 8'd153) ? 1'b0 : ((opcode == 8'd129) ? 1'b0 : ((opcode == 8'd145) ? 1'b0 : ((opcode == 8'd134) ? 1'b0 : ((opcode == 8'd150) ? 1'b0 : ((opcode == 8'd142) ? 1'b0 : ((opcode == 8'd132) ? 1'b0 : ((opcode == 8'd148) ? 1'b0 : ((opcode == 8'd140) ? 1'b0 : ((opcode == 8'd170) ? 1'b0 : ((opcode == 8'd138) ? 1'b0 : ((opcode == 8'd168) ? 1'b0 : ((opcode == 8'd152) ? 1'b0 : ((opcode == 8'd186) ? 1'b0 : ((opcode == 8'd154) ? 1'b0 : ((opcode == 8'd232) ? 1'b0 : ((opcode == 8'd202) ? 1'b0 : ((opcode == 8'd200) ? 1'b0 : ((opcode == 8'd136) ? 1'b0 : ((opcode == 8'd230) ? 1'b0 : ((opcode == 8'd246) ? 1'b0 : ((opcode == 8'd238) ? 1'b0 : ((opcode == 8'd254) ? 1'b0 : ((opcode == 8'd198) ? 1'b0 : ((opcode == 8'd214) ? 1'b0 : ((opcode == 8'd206) ? 1'b0 : ((opcode == 8'd222) ? 1'b0 : ((opcode == 8'd10) ? 1'b0 : ((opcode == 8'd6) ? 1'b0 : ((opcode == 8'd22) ? 1'b0 : ((opcode == 8'd14) ? 1'b0 : ((opcode == 8'd30) ? 1'b0 : ((opcode == 8'd74) ? 1'b0 : ((opcode == 8'd70) ? 1'b0 : ((opcode == 8'd86) ? 1'b0 : ((opcode == 8'd78) ? 1'b0 : ((opcode == 8'd94) ? 1'b0 : ((opcode == 8'd42) ? 1'b0 : ((opcode == 8'd38) ? 1'b0 : ((opcode == 8'd54) ? 1'b0 : ((opcode == 8'd46) ? 1'b0 : ((opcode == 8'd62) ? 1'b0 : ((opcode == 8'd106) ? 1'b0 : ((opcode == 8'd102) ? 1'b0 : ((opcode == 8'd118) ? 1'b0 : ((opcode == 8'd110) ? 1'b0 : ((opcode == 8'd126) ? 1'b0 : ((opcode == 8'd16) ? 1'b0 : ((opcode == 8'd48) ? 1'b0 : ((opcode == 8'd80) ? 1'b0 : ((opcode == 8'd112) ? 1'b0 : ((opcode == 8'd144) ? 1'b0 : ((opcode == 8'd176) ? 1'b0 : ((opcode == 8'd208) ? 1'b0 : ((opcode == 8'd240) ? 1'b0 : ((opcode == 8'd76) ? 1'b0 : ((opcode == 8'd108) ? 1'b0 : ((opcode == 8'd32) ? 1'b0 : ((opcode == 8'd96) ? 1'b0 : ((opcode == 8'd64) ? 1'b0 : ((opcode == 8'd72) ? 1'b0 : ((opcode == 8'd8) ? 1'b0 : ((opcode == 8'd104) ? 1'b0 : ((opcode == 8'd40) ? 1'b0 : ((opcode == 8'd24) ? 1'b0 : ((opcode == 8'd56) ? 1'b0 : ((opcode == 8'd88) ? 1'b0 : ((opcode == 8'd120) ? 1'b0 : ((opcode == 8'd184) ? 1'b0 : ((opcode == 8'd216) ? 1'b0 : ((opcode == 8'd248) ? 1'b0 : ((opcode == 8'd234) ? 1'b0 : ((opcode == 8'd0) ? 1'b0 : 1'b1)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

endmodule