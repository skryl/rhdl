module xnor_gate(
  input a0,
  input a1,
  output y
);

  assign y = ~(a0 ^ a1);

endmodule