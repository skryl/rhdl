module apple2_cpu6502(
  input clk,
  input enable,
  input reset,
  input nmi_n,
  input irq_n,
  input so_n,
  input [7:0] di,
  output [7:0] do_out,
  output [15:0] addr,
  output we,
  output [7:0] debug_opcode,
  output [15:0] debug_pc,
  output [7:0] debug_a,
  output [7:0] debug_x,
  output [7:0] debug_y,
  output [7:0] debug_s,
  output [7:0] debug_p,
  output debug_second_byte,
  output debug_cycle2,
  output [15:0] debug_addr_c2,
  output [47:0] debug_opc_info
);

  reg [4:0] cpu_state;
  reg [7:0] opcode;
  reg [47:0] opc_info;
  reg [7:0] t_reg;
  reg [15:0] pc_reg;
  reg [15:0] addr_reg;
  reg [7:0] a_reg;
  reg [7:0] x_reg;
  reg [7:0] y_reg;
  reg [7:0] s_reg;
  reg flag_c;
  reg flag_z;
  reg flag_i;
  reg flag_d;
  reg flag_v;
  reg flag_n;
  reg irq_active;
  reg nmi_reg;
  reg nmi_edge;
  reg irq_reg;
  reg so_reg;
  reg process_irq;
  reg we_reg;
  reg [7:0] do_reg;
  reg [8:0] index_out;
  reg update_regs;
  wire [4:0] next_state;
  wire [7:0] alu_input;
  wire [7:0] alu_cmp_input;
  wire [7:0] alu_rmw_out;
  wire [7:0] alu_reg_out;
  wire alu_c;
  wire alu_z;
  wire alu_v;
  wire alu_n;
  reg [47:0] opcode_rom [0:255];

  initial begin
    cpu_state = 5'd1;
    opcode = 8'd76;
    opc_info = 48'd66560;
    t_reg = 8'd0;
    pc_reg = 16'd0;
    addr_reg = 16'd65532;
    a_reg = 8'd0;
    x_reg = 8'd0;
    y_reg = 8'd0;
    s_reg = 8'd253;
    flag_c = 1'b0;
    flag_z = 1'b0;
    flag_i = 1'b1;
    flag_d = 1'b0;
    flag_v = 1'b0;
    flag_n = 1'b0;
    irq_active = 1'b0;
    nmi_reg = 1'b1;
    nmi_edge = 1'b1;
    irq_reg = 1'b1;
    so_reg = 1'b1;
    process_irq = 1'b0;
    we_reg = 1'b0;
    do_reg = 8'd0;
  end

  assign addr = addr_reg;
  assign we = we_reg;
  assign do_out = do_reg;
  assign debug_opcode = opcode;
  assign debug_pc = pc_reg;
  assign debug_a = a_reg;
  assign debug_x = x_reg;
  assign debug_y = y_reg;
  assign debug_s = s_reg;
  assign debug_cycle2 = (cpu_state == 5'd1);
  assign debug_second_byte = opc_info[10];
  assign debug_addr_c2 = ((opc_info[10] ? (addr_reg + 16'd1) : addr_reg) & 17'd65535);
  assign debug_opc_info = opc_info;
  assign alu_input = (opc_info[33] ? 8'd0 : (opc_info[31] ? ((opc_info[30] ? ((opc_info[29] ? ((opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255))) & y_reg) : (opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)))) & s_reg) : (opc_info[29] ? ((opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255))) & y_reg) : (opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255))))) & ((enable & (((((cpu_state == 5'd1) | (((cpu_state == 5'd13) | (cpu_state == 5'd14)) & opc_info[20])) | (cpu_state == 5'd4)) | (cpu_state == 5'd8)) | (cpu_state == 5'd9))) ? di : t_reg)) : (opc_info[30] ? ((opc_info[29] ? ((opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255))) & y_reg) : (opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)))) & s_reg) : (opc_info[29] ? ((opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255))) & y_reg) : (opc_info[28] ? ((opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)) & x_reg) : (opc_info[27] ? ((opc_info[26] ? (8'd255 & a_reg) : 8'd255) & (a_reg | 8'd238)) : (opc_info[26] ? (8'd255 & a_reg) : 8'd255)))))));
  assign alu_cmp_input = (opc_info[43] ? ((opc_info[42] ? ((opc_info[41] ? (8'd255 & a_reg) : 8'd255) & x_reg) : (opc_info[41] ? (8'd255 & a_reg) : 8'd255)) & y_reg) : (opc_info[42] ? ((opc_info[41] ? (8'd255 & a_reg) : 8'd255) & x_reg) : (opc_info[41] ? (8'd255 & a_reg) : 8'd255)));
  assign debug_p = {flag_n, flag_v, 1'b1, 1'b0, flag_d, flag_i, flag_z, flag_c};
  assign alu_rmw_out = ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))));
  assign alu_reg_out = ((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))))))));
  assign alu_z = ((opc_info[37:34] == 4'd4) ? ((((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))) >> 1) & 1'b1) : ((((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))))))))) == 8'd0) ? 1'b1 : 1'b0));
  assign alu_n = (((opc_info[37:34] == 4'd5) | (opc_info[37:34] == 4'd4)) ? ((((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))) >> 7) & 1'b1) : ((((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))))))))) >> 7) & 1'b1));
  assign alu_c = ((opc_info[40:38] == 3'd2) ? (((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) >> 8) & 1'b1) : ((opc_info[40:38] == 3'd3) ? (((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) >> 8) & 1'b1) : ((opc_info[40:38] == 3'd1) ? (((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) >> 8) & 1'b1) : ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))))));
  assign alu_v = ((opc_info[40:38] == 3'd2) ? ((a_reg[7] ^ ((((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))))))))) >> 7) & 1'b1)) & (((((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))) >> 7) & 1'b1) ^ ((((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))))))))) >> 7) & 1'b1))) : ((opc_info[40:38] == 3'd3) ? ((a_reg[7] ^ ((((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))))))))) >> 7) & 1'b1)) & (~((((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))) >> 7) & 1'b1) ^ ((((opc_info[40:38] == 3'd2) ? ((({1'b0, a_reg} + {1'b0, ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd3) ? ((({1'b0, a_reg} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, {8'd0, ((((((opc_info[37:34] == 4'd4) | (opc_info[37:34] == 4'd8)) | (opc_info[37:34] == 4'd9)) | (opc_info[37:34] == 4'd10)) | (opc_info[37:34] == 4'd11)) ? ((opc_info[37:34] == 4'd4) ? alu_input[0] : ((opc_info[37:34] == 4'd8) ? alu_input[0] : ((opc_info[37:34] == 4'd9) ? alu_input[0] : ((opc_info[37:34] == 4'd10) ? alu_input[7] : ((opc_info[37:34] == 4'd11) ? alu_input[7] : ((opc_info[37:34] == 4'd15) ? (alu_input[7] & a_reg[7]) : flag_c)))))) : flag_c)}}) & 8'd255) : ((opc_info[40:38] == 3'd1) ? ((({1'b0, alu_cmp_input} + {1'b0, ~((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))}) + {{1{1'b0}}, 9'd1}) & 8'd255) : ((opc_info[40:38] == 3'd4) ? (a_reg & ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd5) ? (a_reg | ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[40:38] == 3'd6) ? (a_reg ^ ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input))))))))))) : ((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))))))))) >> 7) & 1'b1))) : ((opc_info[37:34] == 4'd5) ? ((((opc_info[37:34] == 4'd0) ? alu_input : ((opc_info[37:34] == 4'd1) ? {flag_n, flag_v, 1'b1, ~irq_active, flag_d, flag_i, flag_z, flag_c} : ((opc_info[37:34] == 4'd2) ? ((alu_input + 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd3) ? ((alu_input - 8'd1) & 8'd255) : ((opc_info[37:34] == 4'd4) ? alu_input : ((opc_info[37:34] == 4'd5) ? alu_input : ((opc_info[37:34] == 4'd8) ? {1'b0, alu_input[7:1]} : ((opc_info[37:34] == 4'd9) ? {flag_c, alu_input[7:1]} : ((opc_info[37:34] == 4'd10) ? {alu_input[6:0], 1'b0} : ((opc_info[37:34] == 4'd11) ? {alu_input[6:0], flag_c} : alu_input)))))))))) >> 6) & 1'b1) : alu_input[6])));
  assign next_state = ((cpu_state == 5'd18) ? 5'd0 : ((cpu_state == 5'd17) ? (opc_info[23] ? 5'd18 : 5'd0) : ((cpu_state == 5'd16) ? 5'd8 : ((cpu_state == 5'd15) ? ((~opc_info[15] | opc_info[20]) ? 5'd17 : (opc_info[14] ? 5'd16 : 5'd8)) : ((cpu_state == 5'd14) ? (opc_info[24] ? 5'd8 : ((~opc_info[15] & opc_info[20]) ? 5'd17 : 5'd15)) : ((cpu_state == 5'd13) ? (opc_info[14] ? 5'd14 : 5'd8) : ((cpu_state == 5'd12) ? 5'd0 : ((cpu_state == 5'd11) ? 5'd12 : ((cpu_state == 5'd10) ? 5'd12 : ((cpu_state == 5'd9) ? (opc_info[22] ? 5'd10 : 5'd0) : ((cpu_state == 5'd8) ? (opc_info[16] ? 5'd17 : ((opc_info[17] ? (((({1'b0, t_reg} + {1'b0, pc_reg[7:0]}) >> 8) & 1'b1) ^ t_reg[7]) : ((({1'b0, t_reg} + {1'b0, (opc_info[18] ? x_reg : (opc_info[19] ? y_reg : 8'd0))}) >> 8) & 1'b1)) ? 5'd9 : (opc_info[22] ? ((opc_info[18] | opc_info[19]) ? 5'd9 : 5'd10) : 5'd0))) : ((cpu_state == 5'd7) ? (opc_info[12] ? 5'd9 : 5'd0) : ((cpu_state == 5'd6) ? 5'd0 : ((cpu_state == 5'd5) ? ((opc_info[17] ? (((({1'b0, t_reg} + {1'b0, pc_reg[7:0]}) >> 8) & 1'b1) ^ t_reg[7]) : ((({1'b0, t_reg} + {1'b0, (opc_info[18] ? x_reg : (opc_info[19] ? y_reg : 8'd0))}) >> 8) & 1'b1)) ? 5'd6 : 5'd0) : ((cpu_state == 5'd4) ? 5'd2 : ((cpu_state == 5'd3) ? 5'd4 : ((cpu_state == 5'd2) ? (((opc_info[13] & opc_info[18]) & opc_info[21]) ? 5'd12 : (((opc_info[13] & opc_info[18]) & ~opc_info[21]) ? 5'd9 : ((opc_info[21] & (opc_info[18] | opc_info[19])) ? 5'd11 : ((opc_info[21] & ~(opc_info[18] | opc_info[19])) ? 5'd12 : 5'd8)))) : ((cpu_state == 5'd1) ? ((opc_info[17] & ((opcode[7:6] == 2'd0) ? (flag_n == opcode[5]) : ((opcode[7:6] == 2'd1) ? (flag_v == opcode[5]) : ((opcode[7:6] == 2'd2) ? (flag_c == opcode[5]) : (flag_z == opcode[5]))))) ? 5'd5 : (opc_info[20] ? 5'd13 : ((opc_info[14] & opc_info[15]) ? 5'd14 : ((opc_info[14] & ~opc_info[15]) ? 5'd13 : ((~opc_info[14] & opc_info[15]) ? 5'd12 : (opc_info[11] ? 5'd2 : ((opc_info[13] & opc_info[18]) ? 5'd3 : ((opc_info[13] & ~opc_info[18]) ? 5'd4 : (((opc_info[12] & opc_info[21]) & (opc_info[18] | opc_info[19])) ? 5'd11 : (((opc_info[12] & opc_info[21]) & ~(opc_info[18] | opc_info[19])) ? 5'd12 : (((opc_info[12] & ~opc_info[21]) & (opc_info[18] | opc_info[19])) ? 5'd7 : (((opc_info[12] & ~opc_info[21]) & ~(opc_info[18] | opc_info[19])) ? 5'd9 : (opc_info[16] ? 5'd17 : 5'd0))))))))))))) : ((cpu_state == 5'd0) ? 5'd1 : 5'd0)))))))))))))))))));

  always @(posedge clk) begin
  if (reset) begin
    cpu_state <= 5'd1;
    opcode <= 8'd76;
    opc_info <= 48'd66560;
    t_reg <= 8'd0;
    pc_reg <= 16'd0;
    addr_reg <= 16'd65532;
    a_reg <= 8'd0;
    x_reg <= 8'd0;
    y_reg <= 8'd0;
    s_reg <= 8'd253;
    flag_c <= 1'b0;
    flag_z <= 1'b0;
    flag_i <= 1'b1;
    flag_d <= 1'b0;
    flag_v <= 1'b0;
    flag_n <= 1'b0;
    irq_active <= 1'b0;
    nmi_reg <= 1'b1;
    nmi_edge <= 1'b1;
    irq_reg <= 1'b1;
    so_reg <= 1'b1;
    process_irq <= 1'b0;
    we_reg <= 1'b0;
    do_reg <= 8'd0;
  end
  else begin
    cpu_state <= (enable ? next_state : cpu_state);
    opcode <= ((enable & (cpu_state == 5'd0)) ? (process_irq ? 8'd0 : di) : opcode);
    opc_info <= ((enable & (cpu_state == 5'd0)) ? opcode_rom[(process_irq ? 8'd0 : di)] : opc_info);
    irq_reg <= ((enable & ~((next_state == 5'd5) | (next_state == 5'd0))) ? irq_n : irq_reg);
    nmi_edge <= ((enable & ~((next_state == 5'd5) | (next_state == 5'd0))) ? nmi_n : nmi_edge);
    nmi_reg <= ((enable & (cpu_state == 5'd16)) ? 1'b1 : (((enable & ~((next_state == 5'd5) | (next_state == 5'd0))) & (nmi_edge & ~nmi_n)) ? 1'b0 : nmi_reg));
    process_irq <= (enable ? ~((nmi_reg & (irq_reg | flag_i)) | opc_info[25]) : process_irq);
    irq_active <= ((enable & (cpu_state == 5'd0)) ? (process_irq ? 1'b1 : 1'b0) : irq_active);
    t_reg <= ((enable & (((((cpu_state == 5'd1) | (((cpu_state == 5'd13) | (cpu_state == 5'd14)) & opc_info[20])) | (cpu_state == 5'd4)) | (cpu_state == 5'd8)) | (cpu_state == 5'd9))) ? di : t_reg);
    update_regs <= (opc_info[24] ? (cpu_state == 5'd8) : (next_state == 5'd0));
    a_reg <= (((opc_info[0] & update_regs) & enable) ? alu_reg_out : a_reg);
    x_reg <= (((opc_info[1] & update_regs) & enable) ? alu_reg_out : x_reg);
    y_reg <= (((opc_info[2] & update_regs) & enable) ? alu_reg_out : y_reg);
    s_reg <= (((opc_info[3] & update_regs) & enable) ? alu_reg_out : ((enable & (((((((next_state == 5'd13) & (opc_info[20] | opc_info[15])) | (next_state == 5'd14)) | (next_state == 5'd15)) | (next_state == 5'd16)) | ((next_state == 5'd8) & opc_info[24])) | ((next_state == 5'd12) & opc_info[15]))) ? (opc_info[20] ? ((s_reg + 8'd1) & 8'd255) : ((s_reg - 8'd1) & 8'd255)) : s_reg));
    flag_c <= (((opc_info[9] & update_regs) & enable) ? alu_c : flag_c);
    flag_z <= (((opc_info[8] & update_regs) & enable) ? alu_z : flag_z);
    flag_i <= (((opc_info[7] & update_regs) & enable) ? alu_input[2] : flag_i);
    flag_d <= (((opc_info[6] & update_regs) & enable) ? alu_input[3] : flag_d);
    flag_v <= (((opc_info[5] & update_regs) & enable) ? alu_v : ((enable & (so_reg & ~so_n)) ? 1'b1 : flag_v));
    so_reg <= (enable ? so_n : so_reg);
    flag_n <= (((opc_info[4] & update_regs) & enable) ? alu_n : flag_n);
    pc_reg <= (enable ? ((cpu_state == 5'd0) ? addr_reg : ((((cpu_state == 5'd1) & ~irq_active) & opc_info[10]) ? ((addr_reg + 16'd1) & 16'd65535) : ((((cpu_state == 5'd1) & ~irq_active) & ~opc_info[10]) ? addr_reg : (((cpu_state == 5'd2) & opc_info[11]) ? ((addr_reg + 16'd1) & 16'd65535) : pc_reg)))) : pc_reg);
    we_reg <= (enable ? ((((((next_state == 5'd13) & ~opc_info[20]) & (~opc_info[14] | opc_info[15])) | ((((next_state == 5'd14) | (next_state == 5'd15)) | (next_state == 5'd16)) & ~opc_info[20])) | (next_state == 5'd10)) | (next_state == 5'd12)) : we_reg);
    do_reg <= (enable ? ((next_state == 5'd14) ? ((opc_info[25] & ~irq_active) ? ((((addr_reg + 16'd1) & 16'd65535) >> 8) & 8'd255) : pc_reg[15:8]) : ((next_state == 5'd15) ? pc_reg[7:0] : ((next_state == 5'd10) ? di : (opc_info[32] ? (alu_rmw_out & ((addr_reg[15:8] + 8'd1) & 8'd255)) : alu_rmw_out)))) : do_reg);
    index_out <= (opc_info[17] ? ({1'b0, t_reg} + {1'b0, pc_reg[7:0]}) : ({1'b0, t_reg} + {1'b0, (opc_info[18] ? x_reg : (opc_info[19] ? y_reg : 8'd0))}));
    addr_reg <= (enable ? ((cpu_state == 5'd1) ? ((opc_info[14] | opc_info[15]) ? {8'd1, s_reg} : (opc_info[11] ? ((addr_reg + 16'd1) & 16'd65535) : ((opc_info[12] | opc_info[13]) ? {8'd0, di} : (opc_info[10] ? ((addr_reg + 16'd1) & 16'd65535) : addr_reg)))) : ((cpu_state == 5'd2) ? ((opc_info[13] & opc_info[18]) ? {di, t_reg} : ((opc_info[18] | opc_info[19]) ? {di, ((t_reg + (opc_info[18] ? x_reg : (opc_info[19] ? y_reg : 8'd0))) & 8'd255)} : {di, t_reg})) : ((cpu_state == 5'd3) ? {8'd0, index_out[7:0]} : ((cpu_state == 5'd4) ? {addr_reg[15:8], ((addr_reg[7:0] + 8'd1) & 8'd255)} : ((cpu_state == 5'd5) ? ((pc_reg + (t_reg[7] ? {8'd255, t_reg} : {8'd0, t_reg})) & 16'd65535) : ((cpu_state == 5'd6) ? (t_reg[7] ? {((pc_reg[15:8] - 8'd1) & 8'd255), (((pc_reg + (t_reg[7] ? {8'd255, t_reg} : {8'd0, t_reg})) & 16'd65535) & 8'd255)} : {((pc_reg[15:8] + 8'd1) & 8'd255), (((pc_reg + (t_reg[7] ? {8'd255, t_reg} : {8'd0, t_reg})) & 16'd65535) & 8'd255)}) : ((cpu_state == 5'd7) ? {8'd0, ((t_reg + (opc_info[18] ? x_reg : (opc_info[19] ? y_reg : 8'd0))) & 8'd255)} : ((cpu_state == 5'd8) ? (opc_info[16] ? {addr_reg[15:8], ((addr_reg[7:0] + 8'd1) & 8'd255)} : (index_out[8] ? {((addr_reg[15:8] + 8'd1) & 8'd255), addr_reg[7:0]} : (opc_info[22] ? addr_reg : pc_reg))) : ((cpu_state == 5'd9) ? (opc_info[22] ? addr_reg : pc_reg) : ((cpu_state == 5'd10) ? addr_reg : ((cpu_state == 5'd11) ? (opc_info[12] ? {8'd0, ((t_reg + (opc_info[18] ? x_reg : (opc_info[19] ? y_reg : 8'd0))) & 8'd255)} : (index_out[8] ? {((addr_reg[15:8] + 8'd1) & 8'd255), addr_reg[7:0]} : addr_reg)) : ((cpu_state == 5'd12) ? pc_reg : (((cpu_state == 5'd13) | (cpu_state == 5'd14)) ? {8'd1, s_reg} : ((cpu_state == 5'd15) ? (opc_info[16] ? pc_reg : {8'd1, s_reg}) : ((cpu_state == 5'd16) ? (nmi_reg ? 16'd65534 : 16'd65530) : ((cpu_state == 5'd17) ? {di, t_reg} : ((addr_reg + 16'd1) & 16'd65535))))))))))))))))) : addr_reg);
  end
  end

endmodule