module alu #(
  parameter width = 8
) (
  input [7:0] a,
  input [7:0] b,
  input [3:0] op,
  input cin,
  output [7:0] result,
  output cout,
  output zero,
  output negative,
  output overflow
);

  assign result = ((op == 4'd0) ? (((a + b) + {{8{1'b0}}, cin}) & 8'd255) : ((op == 4'd1) ? (((a - b) - {{7{1'b0}}, cin}) & 8'd255) : ((op == 4'd2) ? (a & b) : ((op == 4'd3) ? (a | b) : ((op == 4'd4) ? (a ^ b) : ((op == 4'd5) ? ~a : ((op == 4'd6) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[6:0], 1'b0} : ((b[2:0] == 3'd2) ? {a[5:0], 2'd0} : ((b[2:0] == 3'd3) ? {a[4:0], 3'd0} : ((b[2:0] == 3'd4) ? {a[3:0], 4'd0} : ((b[2:0] == 3'd5) ? {a[2:0], 5'd0} : ((b[2:0] == 3'd6) ? {a[1:0], 6'd0} : ((b[2:0] == 3'd7) ? {a[0], 7'd0} : a)))))))) : ((op == 4'd7) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {1'b0, a[7:1]} : ((b[2:0] == 3'd2) ? {2'd0, a[7:2]} : ((b[2:0] == 3'd3) ? {3'd0, a[7:3]} : ((b[2:0] == 3'd4) ? {4'd0, a[7:4]} : ((b[2:0] == 3'd5) ? {5'd0, a[7:5]} : ((b[2:0] == 3'd6) ? {6'd0, a[7:6]} : ((b[2:0] == 3'd7) ? {7'd0, a[7]} : a)))))))) : ((op == 4'd8) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[7], a[7:1]} : ((b[2:0] == 3'd2) ? {{a[7], a[7]}, a[7:2]} : ((b[2:0] == 3'd3) ? {{a[7], a[7], a[7]}, a[7:3]} : ((b[2:0] == 3'd4) ? {{a[7], a[7], a[7], a[7]}, a[7:4]} : ((b[2:0] == 3'd5) ? {{a[7], a[7], a[7], a[7], a[7]}, a[7:5]} : ((b[2:0] == 3'd6) ? {{a[7], a[7], a[7], a[7], a[7], a[7]}, a[7:6]} : ((b[2:0] == 3'd7) ? {{a[7], a[7], a[7], a[7], a[7], a[7], a[7]}, a[7]} : a)))))))) : ((op == 4'd9) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[6:0], a[7]} : ((b[2:0] == 3'd2) ? {a[5:0], a[7:6]} : ((b[2:0] == 3'd3) ? {a[4:0], a[7:5]} : ((b[2:0] == 3'd4) ? {a[3:0], a[7:4]} : ((b[2:0] == 3'd5) ? {a[2:0], a[7:3]} : ((b[2:0] == 3'd6) ? {a[1:0], a[7:2]} : ((b[2:0] == 3'd7) ? {a[0], a[7:1]} : a)))))))) : ((op == 4'd10) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[0], a[7:1]} : ((b[2:0] == 3'd2) ? {a[1:0], a[7:2]} : ((b[2:0] == 3'd3) ? {a[2:0], a[7:3]} : ((b[2:0] == 3'd4) ? {a[3:0], a[7:4]} : ((b[2:0] == 3'd5) ? {a[4:0], a[7:5]} : ((b[2:0] == 3'd6) ? {a[5:0], a[7:6]} : ((b[2:0] == 3'd7) ? {a[6:0], a[7]} : a)))))))) : ((op == 4'd11) ? ((a * b) & 8'd255) : ((op == 4'd12) ? (a / b) : ((op == 4'd13) ? (a % b) : ((op == 4'd14) ? ((a + 8'd1) & 8'd255) : ((op == 4'd15) ? ((a - 8'd1) & 8'd255) : (((a + b) + {{8{1'b0}}, cin}) & 8'd255)))))))))))))))));
  assign cout = ((op == 4'd0) ? ((((a + b) + {{8{1'b0}}, cin}) >> 8) & 1'b1) : ((op == 4'd1) ? ((a < ((b + {{7{1'b0}}, cin}) & 9'd255)) ? 1'b1 : 1'b0) : ((op == 4'd2) ? 1'b0 : ((op == 4'd3) ? 1'b0 : ((op == 4'd4) ? 1'b0 : ((op == 4'd5) ? 1'b0 : ((op == 4'd6) ? a[7] : ((op == 4'd7) ? a[0] : ((op == 4'd8) ? a[0] : ((op == 4'd9) ? a[7] : ((op == 4'd10) ? a[0] : ((op == 4'd11) ? (((((a * b) >> 8) & 8'd255) != 8'd0) ? 1'b1 : 1'b0) : ((op == 4'd12) ? ((b == 8'd0) ? 1'b1 : 1'b0) : ((op == 4'd13) ? ((b == 8'd0) ? 1'b1 : 1'b0) : ((op == 4'd14) ? (((a + 8'd1) >> 8) & 1'b1) : ((op == 4'd15) ? ((a == 8'd0) ? 1'b1 : 1'b0) : ((((a + b) + {{8{1'b0}}, cin}) >> 8) & 1'b1)))))))))))))))));
  assign overflow = ((op == 4'd0) ? ((a[7] == b[7]) & ((((((a + b) + {{8{1'b0}}, cin}) & 8'd255) >> 7) & 1'b1) != a[7])) : ((op == 4'd1) ? ((a[7] != b[7]) & ((((((a - b) - {{7{1'b0}}, cin}) & 8'd255) >> 7) & 1'b1) != a[7])) : ((op == 4'd2) ? 1'b0 : ((op == 4'd3) ? 1'b0 : ((op == 4'd4) ? 1'b0 : ((op == 4'd5) ? 1'b0 : ((op == 4'd6) ? 1'b0 : ((op == 4'd7) ? 1'b0 : ((op == 4'd8) ? 1'b0 : ((op == 4'd9) ? 1'b0 : ((op == 4'd10) ? 1'b0 : ((op == 4'd11) ? 1'b0 : ((op == 4'd12) ? 1'b0 : ((op == 4'd13) ? 1'b0 : ((op == 4'd14) ? ((a == 8'd127) ? 1'b1 : 1'b0) : ((op == 4'd15) ? ((a == 8'd128) ? 1'b1 : 1'b0) : ((a[7] == b[7]) & ((((((a + b) + {{8{1'b0}}, cin}) & 8'd255) >> 7) & 1'b1) != a[7]))))))))))))))))));
  assign zero = ((((op == 4'd0) ? (((a + b) + {{8{1'b0}}, cin}) & 8'd255) : ((op == 4'd1) ? (((a - b) - {{7{1'b0}}, cin}) & 8'd255) : ((op == 4'd2) ? (a & b) : ((op == 4'd3) ? (a | b) : ((op == 4'd4) ? (a ^ b) : ((op == 4'd5) ? ~a : ((op == 4'd6) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[6:0], 1'b0} : ((b[2:0] == 3'd2) ? {a[5:0], 2'd0} : ((b[2:0] == 3'd3) ? {a[4:0], 3'd0} : ((b[2:0] == 3'd4) ? {a[3:0], 4'd0} : ((b[2:0] == 3'd5) ? {a[2:0], 5'd0} : ((b[2:0] == 3'd6) ? {a[1:0], 6'd0} : ((b[2:0] == 3'd7) ? {a[0], 7'd0} : a)))))))) : ((op == 4'd7) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {1'b0, a[7:1]} : ((b[2:0] == 3'd2) ? {2'd0, a[7:2]} : ((b[2:0] == 3'd3) ? {3'd0, a[7:3]} : ((b[2:0] == 3'd4) ? {4'd0, a[7:4]} : ((b[2:0] == 3'd5) ? {5'd0, a[7:5]} : ((b[2:0] == 3'd6) ? {6'd0, a[7:6]} : ((b[2:0] == 3'd7) ? {7'd0, a[7]} : a)))))))) : ((op == 4'd8) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[7], a[7:1]} : ((b[2:0] == 3'd2) ? {{a[7], a[7]}, a[7:2]} : ((b[2:0] == 3'd3) ? {{a[7], a[7], a[7]}, a[7:3]} : ((b[2:0] == 3'd4) ? {{a[7], a[7], a[7], a[7]}, a[7:4]} : ((b[2:0] == 3'd5) ? {{a[7], a[7], a[7], a[7], a[7]}, a[7:5]} : ((b[2:0] == 3'd6) ? {{a[7], a[7], a[7], a[7], a[7], a[7]}, a[7:6]} : ((b[2:0] == 3'd7) ? {{a[7], a[7], a[7], a[7], a[7], a[7], a[7]}, a[7]} : a)))))))) : ((op == 4'd9) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[6:0], a[7]} : ((b[2:0] == 3'd2) ? {a[5:0], a[7:6]} : ((b[2:0] == 3'd3) ? {a[4:0], a[7:5]} : ((b[2:0] == 3'd4) ? {a[3:0], a[7:4]} : ((b[2:0] == 3'd5) ? {a[2:0], a[7:3]} : ((b[2:0] == 3'd6) ? {a[1:0], a[7:2]} : ((b[2:0] == 3'd7) ? {a[0], a[7:1]} : a)))))))) : ((op == 4'd10) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[0], a[7:1]} : ((b[2:0] == 3'd2) ? {a[1:0], a[7:2]} : ((b[2:0] == 3'd3) ? {a[2:0], a[7:3]} : ((b[2:0] == 3'd4) ? {a[3:0], a[7:4]} : ((b[2:0] == 3'd5) ? {a[4:0], a[7:5]} : ((b[2:0] == 3'd6) ? {a[5:0], a[7:6]} : ((b[2:0] == 3'd7) ? {a[6:0], a[7]} : a)))))))) : ((op == 4'd11) ? ((a * b) & 8'd255) : ((op == 4'd12) ? (a / b) : ((op == 4'd13) ? (a % b) : ((op == 4'd14) ? ((a + 8'd1) & 8'd255) : ((op == 4'd15) ? ((a - 8'd1) & 8'd255) : (((a + b) + {{8{1'b0}}, cin}) & 8'd255))))))))))))))))) == 8'd0) ? 1'b1 : 1'b0);
  assign negative = ((((op == 4'd0) ? (((a + b) + {{8{1'b0}}, cin}) & 8'd255) : ((op == 4'd1) ? (((a - b) - {{7{1'b0}}, cin}) & 8'd255) : ((op == 4'd2) ? (a & b) : ((op == 4'd3) ? (a | b) : ((op == 4'd4) ? (a ^ b) : ((op == 4'd5) ? ~a : ((op == 4'd6) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[6:0], 1'b0} : ((b[2:0] == 3'd2) ? {a[5:0], 2'd0} : ((b[2:0] == 3'd3) ? {a[4:0], 3'd0} : ((b[2:0] == 3'd4) ? {a[3:0], 4'd0} : ((b[2:0] == 3'd5) ? {a[2:0], 5'd0} : ((b[2:0] == 3'd6) ? {a[1:0], 6'd0} : ((b[2:0] == 3'd7) ? {a[0], 7'd0} : a)))))))) : ((op == 4'd7) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {1'b0, a[7:1]} : ((b[2:0] == 3'd2) ? {2'd0, a[7:2]} : ((b[2:0] == 3'd3) ? {3'd0, a[7:3]} : ((b[2:0] == 3'd4) ? {4'd0, a[7:4]} : ((b[2:0] == 3'd5) ? {5'd0, a[7:5]} : ((b[2:0] == 3'd6) ? {6'd0, a[7:6]} : ((b[2:0] == 3'd7) ? {7'd0, a[7]} : a)))))))) : ((op == 4'd8) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[7], a[7:1]} : ((b[2:0] == 3'd2) ? {{a[7], a[7]}, a[7:2]} : ((b[2:0] == 3'd3) ? {{a[7], a[7], a[7]}, a[7:3]} : ((b[2:0] == 3'd4) ? {{a[7], a[7], a[7], a[7]}, a[7:4]} : ((b[2:0] == 3'd5) ? {{a[7], a[7], a[7], a[7], a[7]}, a[7:5]} : ((b[2:0] == 3'd6) ? {{a[7], a[7], a[7], a[7], a[7], a[7]}, a[7:6]} : ((b[2:0] == 3'd7) ? {{a[7], a[7], a[7], a[7], a[7], a[7], a[7]}, a[7]} : a)))))))) : ((op == 4'd9) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[6:0], a[7]} : ((b[2:0] == 3'd2) ? {a[5:0], a[7:6]} : ((b[2:0] == 3'd3) ? {a[4:0], a[7:5]} : ((b[2:0] == 3'd4) ? {a[3:0], a[7:4]} : ((b[2:0] == 3'd5) ? {a[2:0], a[7:3]} : ((b[2:0] == 3'd6) ? {a[1:0], a[7:2]} : ((b[2:0] == 3'd7) ? {a[0], a[7:1]} : a)))))))) : ((op == 4'd10) ? ((b[2:0] == 3'd0) ? a : ((b[2:0] == 3'd1) ? {a[0], a[7:1]} : ((b[2:0] == 3'd2) ? {a[1:0], a[7:2]} : ((b[2:0] == 3'd3) ? {a[2:0], a[7:3]} : ((b[2:0] == 3'd4) ? {a[3:0], a[7:4]} : ((b[2:0] == 3'd5) ? {a[4:0], a[7:5]} : ((b[2:0] == 3'd6) ? {a[5:0], a[7:6]} : ((b[2:0] == 3'd7) ? {a[6:0], a[7]} : a)))))))) : ((op == 4'd11) ? ((a * b) & 8'd255) : ((op == 4'd12) ? (a / b) : ((op == 4'd13) ? (a % b) : ((op == 4'd14) ? ((a + 8'd1) & 8'd255) : ((op == 4'd15) ? ((a - 8'd1) & 8'd255) : (((a + b) + {{8{1'b0}}, cin}) & 8'd255))))))))))))))))) >> 7) & 1'b1);

endmodule