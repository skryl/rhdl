library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bitwise_not is
  port(
    a : in std_logic_vector(7 downto 0);
    y : out std_logic_vector(7 downto 0)
  );
end bitwise_not;

architecture rtl of bitwise_not is
begin
  y <= not a;
end rtl;