module memory_address_register
  (
    input clk,
    input reset,
    input load,
    input increment,
    input [7:0] data_in,
    output [7:0] data_out,
    input clk,
    input reset,
    input [7:0] a,
    input [7:0] b,
    input [3:0] op,
    output [7:0] result,
    output zero_flag,
    input clk,
    input reset,
    input [7:0] address,
    input [7:0] data_in,
    input write_enable,
    output [7:0] data_out,
    input clk,
    input reset,
    input [7:0] data_in,
    input load,
    output [7:0] data_out
  );


endmodule